module cla_4bits (
    input   [3 : 0]     p,g             ,
    input               cin             ,
    output  [3 : 0]     s               ,
    output              pout,gout,cout
);

endmodule